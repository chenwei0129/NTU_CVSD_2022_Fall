module XOR_u(
  input clk_i,
  input rst_ni,
  input en_i,
  input u0_i,
  input u1_i,
  input [8:0] select_i,
  input [2:0] select_o_i,
  output reg [255:0]  u_o
);
  
  reg [511:0] u;
  wire [9:0] index = select_i << 1;
  
  reg [255:0] u0_o ;
  //reg [511:0] u0_t ;
  reg [509:0] u0_t ;
  reg [255:0] u1_o ;
  //reg [511:0] u1_t ;
  reg [507:0] u1_t ;
  reg [255:0] u2_o ;
  //reg [511:0] u2_t ;
  reg [503:0] u2_t ;
  reg [255:0] u3_o ;
  //reg [511:0] u3_t ;
  reg [495:0] u3_t ;
  reg [255:0] u4_o ;
  //reg [511:0] u4_t ;
  reg [479:0] u4_t ;
  reg [255:0] u5_o ;
  //reg [511:0] u5_t ;
  reg [447:0] u5_t ;
  reg [255:0] u6_o ;
  //reg [511:0] u6_t ;
  reg [383:0] u6_t ;
  reg [255:0] u7_o ;
  //reg [511:0] u7_t ;
  reg [255:0] u7_t ;
  
  always@(*)begin
    case(select_o_i)
      3'd7   :u_o = u7_o;
      3'd6   :u_o = u6_o;
      3'd5   :u_o = u5_o;
      3'd4   :u_o = u4_o;
      3'd3   :u_o = u3_o;
      3'd2   :u_o = u2_o;
      3'd1   :u_o = u1_o;
      default:u_o = u0_o;
    endcase
  end
  
  integer i;
  always@(posedge clk_i)begin
    if(rst_ni)begin
      for(i=0;i<512;i=i+1)begin
        u[i] <= 1'b0;
      end
    end else if(en_i)begin
      u[index]      <= u0_i;
      u[index+1] <= u1_i;
    end
  end
  
  always@(posedge clk_i)begin
    for(i=0;i<256;i=i+2)begin
      u0_o[i]   <= u0_t[i*2];
      u0_o[i+1] <= u0_t[i*2+1];
    end
  end
  
  always@(posedge clk_i)begin
    for(i=0;i<256;i=i+4)begin
      u1_o[i]   <= u1_t[i*2];
      u1_o[i+1] <= u1_t[i*2+1];
      u1_o[i+2] <= u1_t[i*2+2];
      u1_o[i+3] <= u1_t[i*2+3];
    end
  end
  
  always@(posedge clk_i)begin
    for(i=0;i<256;i=i+8)begin
      u2_o[i]   <= u2_t[i*2];
      u2_o[i+1] <= u2_t[i*2+1];
      u2_o[i+2] <= u2_t[i*2+2];
      u2_o[i+3] <= u2_t[i*2+3];
      u2_o[i+4] <= u2_t[i*2+4];
      u2_o[i+5] <= u2_t[i*2+5];
      u2_o[i+6] <= u2_t[i*2+6];
      u2_o[i+7] <= u2_t[i*2+7];
    end
  end
  
  always@(posedge clk_i)begin
    for(i=0;i<256;i=i+16)begin
      u3_o[i]    <= u3_t[i*2];
      u3_o[i+1]  <= u3_t[i*2+1];
      u3_o[i+2]  <= u3_t[i*2+2];
      u3_o[i+3]  <= u3_t[i*2+3];
      u3_o[i+4]  <= u3_t[i*2+4];
      u3_o[i+5]  <= u3_t[i*2+5];
      u3_o[i+6]  <= u3_t[i*2+6];
      u3_o[i+7]  <= u3_t[i*2+7];
      u3_o[i+8]  <= u3_t[i*2+8];
      u3_o[i+9]  <= u3_t[i*2+9];
      u3_o[i+10] <= u3_t[i*2+10];
      u3_o[i+11] <= u3_t[i*2+11];
      u3_o[i+12] <= u3_t[i*2+12];
      u3_o[i+13] <= u3_t[i*2+13];
      u3_o[i+14] <= u3_t[i*2+14];
      u3_o[i+15] <= u3_t[i*2+15];
    end
  end
  
  always@(posedge clk_i)begin
    for(i=0;i<256;i=i+32)begin
      u4_o[i]    <= u4_t[i*2];
      u4_o[i+1]  <= u4_t[i*2+1];
      u4_o[i+2]  <= u4_t[i*2+2];
      u4_o[i+3]  <= u4_t[i*2+3];
      u4_o[i+4]  <= u4_t[i*2+4];
      u4_o[i+5]  <= u4_t[i*2+5];
      u4_o[i+6]  <= u4_t[i*2+6];
      u4_o[i+7]  <= u4_t[i*2+7];
      u4_o[i+8]  <= u4_t[i*2+8];
      u4_o[i+9]  <= u4_t[i*2+9];
      u4_o[i+10] <= u4_t[i*2+10];
      u4_o[i+11] <= u4_t[i*2+11];
      u4_o[i+12] <= u4_t[i*2+12];
      u4_o[i+13] <= u4_t[i*2+13];
      u4_o[i+14] <= u4_t[i*2+14];
      u4_o[i+15] <= u4_t[i*2+15];
      u4_o[i+16] <= u4_t[i*2+16];
      u4_o[i+17] <= u4_t[i*2+17];
      u4_o[i+18] <= u4_t[i*2+18];
      u4_o[i+19] <= u4_t[i*2+19];
      u4_o[i+20] <= u4_t[i*2+20];
      u4_o[i+21] <= u4_t[i*2+21];
      u4_o[i+22] <= u4_t[i*2+22];
      u4_o[i+23] <= u4_t[i*2+23];
      u4_o[i+24] <= u4_t[i*2+24];
      u4_o[i+25] <= u4_t[i*2+25];
      u4_o[i+26] <= u4_t[i*2+26];
      u4_o[i+27] <= u4_t[i*2+27];
      u4_o[i+28] <= u4_t[i*2+28];
      u4_o[i+29] <= u4_t[i*2+29];
      u4_o[i+30] <= u4_t[i*2+30];
      u4_o[i+31] <= u4_t[i*2+31];
    end
  end
  
  always@(posedge clk_i)begin
    for(i=0;i<256;i=i+64)begin
      u5_o[i]  <= u5_t[i*2];
      u5_o[i+1]  <= u5_t[i*2+1];
      u5_o[i+2]  <= u5_t[i*2+2];
      u5_o[i+3]  <= u5_t[i*2+3];
      u5_o[i+4]  <= u5_t[i*2+4];
      u5_o[i+5]  <= u5_t[i*2+5];
      u5_o[i+6]  <= u5_t[i*2+6];
      u5_o[i+7]  <= u5_t[i*2+7];
      u5_o[i+8]  <= u5_t[i*2+8];
      u5_o[i+9]  <= u5_t[i*2+9];
      u5_o[i+10] <= u5_t[i*2+10];
      u5_o[i+11] <= u5_t[i*2+11];
      u5_o[i+12] <= u5_t[i*2+12];
      u5_o[i+13] <= u5_t[i*2+13];
      u5_o[i+14] <= u5_t[i*2+14];
      u5_o[i+15] <= u5_t[i*2+15];
      u5_o[i+16] <= u5_t[i*2+16];
      u5_o[i+17] <= u5_t[i*2+17];
      u5_o[i+18] <= u5_t[i*2+18];
      u5_o[i+19] <= u5_t[i*2+19];
      u5_o[i+20] <= u5_t[i*2+20];
      u5_o[i+21] <= u5_t[i*2+21];
      u5_o[i+22] <= u5_t[i*2+22];
      u5_o[i+23] <= u5_t[i*2+23];
      u5_o[i+24] <= u5_t[i*2+24];
      u5_o[i+25] <= u5_t[i*2+25];
      u5_o[i+26] <= u5_t[i*2+26];
      u5_o[i+27] <= u5_t[i*2+27];
      u5_o[i+28] <= u5_t[i*2+28];
      u5_o[i+29] <= u5_t[i*2+29];
      u5_o[i+30] <= u5_t[i*2+30];
      u5_o[i+31] <= u5_t[i*2+31];
      u5_o[i+32] <= u5_t[i*2+32];
      u5_o[i+33] <= u5_t[i*2+33];
      u5_o[i+34] <= u5_t[i*2+34];
      u5_o[i+35] <= u5_t[i*2+35];
      u5_o[i+36] <= u5_t[i*2+36];
      u5_o[i+37] <= u5_t[i*2+37];
      u5_o[i+38] <= u5_t[i*2+38];
      u5_o[i+39] <= u5_t[i*2+39];
      u5_o[i+40] <= u5_t[i*2+40];
      u5_o[i+41] <= u5_t[i*2+41];
      u5_o[i+42] <= u5_t[i*2+42];
      u5_o[i+43] <= u5_t[i*2+43];
      u5_o[i+44] <= u5_t[i*2+44];
      u5_o[i+45] <= u5_t[i*2+45];
      u5_o[i+46] <= u5_t[i*2+46];
      u5_o[i+47] <= u5_t[i*2+47];
      u5_o[i+48] <= u5_t[i*2+48];
      u5_o[i+49] <= u5_t[i*2+49];
      u5_o[i+50] <= u5_t[i*2+50];
      u5_o[i+51] <= u5_t[i*2+51];
      u5_o[i+52] <= u5_t[i*2+52];
      u5_o[i+53] <= u5_t[i*2+53];
      u5_o[i+54] <= u5_t[i*2+54];
      u5_o[i+55] <= u5_t[i*2+55];
      u5_o[i+56] <= u5_t[i*2+56];
      u5_o[i+57] <= u5_t[i*2+57];
      u5_o[i+58] <= u5_t[i*2+58];
      u5_o[i+59] <= u5_t[i*2+59];
      u5_o[i+60] <= u5_t[i*2+60];
      u5_o[i+61] <= u5_t[i*2+61];
      u5_o[i+62] <= u5_t[i*2+62];
      u5_o[i+63] <= u5_t[i*2+63];
    end
  end
  
  always@(posedge clk_i)begin
    for(i=0;i<256;i=i+128)begin
      u6_o[i]  <= u6_t[i*2];
      u6_o[i+1]  <= u6_t[i*2+1];
      u6_o[i+2]  <= u6_t[i*2+2];
      u6_o[i+3]  <= u6_t[i*2+3];
      u6_o[i+4]  <= u6_t[i*2+4];
      u6_o[i+5]  <= u6_t[i*2+5];
      u6_o[i+6]  <= u6_t[i*2+6];
      u6_o[i+7]  <= u6_t[i*2+7];
      u6_o[i+8]  <= u6_t[i*2+8];
      u6_o[i+9]  <= u6_t[i*2+9];
      u6_o[i+10] <= u6_t[i*2+10];
      u6_o[i+11] <= u6_t[i*2+11];
      u6_o[i+12] <= u6_t[i*2+12];
      u6_o[i+13] <= u6_t[i*2+13];
      u6_o[i+14] <= u6_t[i*2+14];
      u6_o[i+15] <= u6_t[i*2+15];
      u6_o[i+16] <= u6_t[i*2+16];
      u6_o[i+17] <= u6_t[i*2+17];
      u6_o[i+18] <= u6_t[i*2+18];
      u6_o[i+19] <= u6_t[i*2+19];
      u6_o[i+20] <= u6_t[i*2+20];
      u6_o[i+21] <= u6_t[i*2+21];
      u6_o[i+22] <= u6_t[i*2+22];
      u6_o[i+23] <= u6_t[i*2+23];
      u6_o[i+24] <= u6_t[i*2+24];
      u6_o[i+25] <= u6_t[i*2+25];
      u6_o[i+26] <= u6_t[i*2+26];
      u6_o[i+27] <= u6_t[i*2+27];
      u6_o[i+28] <= u6_t[i*2+28];
      u6_o[i+29] <= u6_t[i*2+29];
      u6_o[i+30] <= u6_t[i*2+30];
      u6_o[i+31] <= u6_t[i*2+31];
      u6_o[i+32] <= u6_t[i*2+32];
      u6_o[i+33] <= u6_t[i*2+33];
      u6_o[i+34] <= u6_t[i*2+34];
      u6_o[i+35] <= u6_t[i*2+35];
      u6_o[i+36] <= u6_t[i*2+36];
      u6_o[i+37] <= u6_t[i*2+37];
      u6_o[i+38] <= u6_t[i*2+38];
      u6_o[i+39] <= u6_t[i*2+39];
      u6_o[i+40] <= u6_t[i*2+40];
      u6_o[i+41] <= u6_t[i*2+41];
      u6_o[i+42] <= u6_t[i*2+42];
      u6_o[i+43] <= u6_t[i*2+43];
      u6_o[i+44] <= u6_t[i*2+44];
      u6_o[i+45] <= u6_t[i*2+45];
      u6_o[i+46] <= u6_t[i*2+46];
      u6_o[i+47] <= u6_t[i*2+47];
      u6_o[i+48] <= u6_t[i*2+48];
      u6_o[i+49] <= u6_t[i*2+49];
      u6_o[i+50] <= u6_t[i*2+50];
      u6_o[i+51] <= u6_t[i*2+51];
      u6_o[i+52] <= u6_t[i*2+52];
      u6_o[i+53] <= u6_t[i*2+53];
      u6_o[i+54] <= u6_t[i*2+54];
      u6_o[i+55] <= u6_t[i*2+55];
      u6_o[i+56] <= u6_t[i*2+56];
      u6_o[i+57] <= u6_t[i*2+57];
      u6_o[i+58] <= u6_t[i*2+58];
      u6_o[i+59] <= u6_t[i*2+59];
      u6_o[i+60] <= u6_t[i*2+60];
      u6_o[i+61] <= u6_t[i*2+61];
      u6_o[i+62] <= u6_t[i*2+62];
      u6_o[i+63] <= u6_t[i*2+63];
      u6_o[i+64] <= u6_t[i*2+64];
      u6_o[i+65] <= u6_t[i*2+65];
      u6_o[i+66] <= u6_t[i*2+66];
      u6_o[i+67] <= u6_t[i*2+67];
      u6_o[i+68] <= u6_t[i*2+68];
      u6_o[i+69] <= u6_t[i*2+69];
      u6_o[i+70] <= u6_t[i*2+70];
      u6_o[i+71] <= u6_t[i*2+71];
      u6_o[i+72] <= u6_t[i*2+72];
      u6_o[i+73] <= u6_t[i*2+73];
      u6_o[i+74] <= u6_t[i*2+74];
      u6_o[i+75] <= u6_t[i*2+75];
      u6_o[i+76] <= u6_t[i*2+76];
      u6_o[i+77] <= u6_t[i*2+77];
      u6_o[i+78] <= u6_t[i*2+78];
      u6_o[i+79] <= u6_t[i*2+79];
      u6_o[i+80] <= u6_t[i*2+80];
      u6_o[i+81] <= u6_t[i*2+81];
      u6_o[i+82] <= u6_t[i*2+82];
      u6_o[i+83] <= u6_t[i*2+83];
      u6_o[i+84] <= u6_t[i*2+84];
      u6_o[i+85] <= u6_t[i*2+85];
      u6_o[i+86] <= u6_t[i*2+86];
      u6_o[i+87] <= u6_t[i*2+87];
      u6_o[i+88] <= u6_t[i*2+88];
      u6_o[i+89] <= u6_t[i*2+89];
      u6_o[i+90] <= u6_t[i*2+90];
      u6_o[i+91] <= u6_t[i*2+91];
      u6_o[i+92] <= u6_t[i*2+92];
      u6_o[i+93] <= u6_t[i*2+93];
      u6_o[i+94] <= u6_t[i*2+94];
      u6_o[i+95] <= u6_t[i*2+95];
      u6_o[i+96] <= u6_t[i*2+96];
      u6_o[i+97] <= u6_t[i*2+97];
      u6_o[i+98] <= u6_t[i*2+98];
      u6_o[i+99] <= u6_t[i*2+99];
      u6_o[i+100] <= u6_t[i*2+100];
      u6_o[i+101] <= u6_t[i*2+101];
      u6_o[i+102] <= u6_t[i*2+102];
      u6_o[i+103] <= u6_t[i*2+103];
      u6_o[i+104] <= u6_t[i*2+104];
      u6_o[i+105] <= u6_t[i*2+105];
      u6_o[i+106] <= u6_t[i*2+106];
      u6_o[i+107] <= u6_t[i*2+107];
      u6_o[i+108] <= u6_t[i*2+108];
      u6_o[i+109] <= u6_t[i*2+109];
      u6_o[i+110] <= u6_t[i*2+110];
      u6_o[i+111] <= u6_t[i*2+111];
      u6_o[i+112] <= u6_t[i*2+112];
      u6_o[i+113] <= u6_t[i*2+113];
      u6_o[i+114] <= u6_t[i*2+114];
      u6_o[i+115] <= u6_t[i*2+115];
      u6_o[i+116] <= u6_t[i*2+116];
      u6_o[i+117] <= u6_t[i*2+117];
      u6_o[i+118] <= u6_t[i*2+118];
      u6_o[i+119] <= u6_t[i*2+119];
      u6_o[i+120] <= u6_t[i*2+120];
      u6_o[i+121] <= u6_t[i*2+121];
      u6_o[i+122] <= u6_t[i*2+122];
      u6_o[i+123] <= u6_t[i*2+123];
      u6_o[i+124] <= u6_t[i*2+124];
      u6_o[i+125] <= u6_t[i*2+125];
      u6_o[i+126] <= u6_t[i*2+126];
      u6_o[i+127] <= u6_t[i*2+127];
    end
  end
  
  always@(posedge clk_i)begin
    u7_o[0]  <= u7_t[0];
    u7_o[1]  <= u7_t[1];
    u7_o[2]  <= u7_t[2];
    u7_o[3]  <= u7_t[3];
    u7_o[4]  <= u7_t[4];
    u7_o[5]  <= u7_t[5];
    u7_o[6]  <= u7_t[6];
    u7_o[7]  <= u7_t[7];
    u7_o[8]  <= u7_t[8];
    u7_o[9]  <= u7_t[9];
    u7_o[10] <= u7_t[10];
    u7_o[11] <= u7_t[11];
    u7_o[12] <= u7_t[12];
    u7_o[13] <= u7_t[13];
    u7_o[14] <= u7_t[14];
    u7_o[15] <= u7_t[15];
    u7_o[16] <= u7_t[16];
    u7_o[17] <= u7_t[17];
    u7_o[18] <= u7_t[18];
    u7_o[19] <= u7_t[19];
    u7_o[20] <= u7_t[20];
    u7_o[21] <= u7_t[21];
    u7_o[22] <= u7_t[22];
    u7_o[23] <= u7_t[23];
    u7_o[24] <= u7_t[24];
    u7_o[25] <= u7_t[25];
    u7_o[26] <= u7_t[26];
    u7_o[27] <= u7_t[27];
    u7_o[28] <= u7_t[28];
    u7_o[29] <= u7_t[29];
    u7_o[30] <= u7_t[30];
    u7_o[31] <= u7_t[31];
    u7_o[32] <= u7_t[32];
    u7_o[33] <= u7_t[33];
    u7_o[34] <= u7_t[34];
    u7_o[35] <= u7_t[35];
    u7_o[36] <= u7_t[36];
    u7_o[37] <= u7_t[37];
    u7_o[38] <= u7_t[38];
    u7_o[39] <= u7_t[39];
    u7_o[40] <= u7_t[40];
    u7_o[41] <= u7_t[41];
    u7_o[42] <= u7_t[42];
    u7_o[43] <= u7_t[43];
    u7_o[44] <= u7_t[44];
    u7_o[45] <= u7_t[45];
    u7_o[46] <= u7_t[46];
    u7_o[47] <= u7_t[47];
    u7_o[48] <= u7_t[48];
    u7_o[49] <= u7_t[49];
    u7_o[50] <= u7_t[50];
    u7_o[51] <= u7_t[51];
    u7_o[52] <= u7_t[52];
    u7_o[53] <= u7_t[53];
    u7_o[54] <= u7_t[54];
    u7_o[55] <= u7_t[55];
    u7_o[56] <= u7_t[56];
    u7_o[57] <= u7_t[57];
    u7_o[58] <= u7_t[58];
    u7_o[59] <= u7_t[59];
    u7_o[60] <= u7_t[60];
    u7_o[61] <= u7_t[61];
    u7_o[62] <= u7_t[62];
    u7_o[63] <= u7_t[63];
    u7_o[64] <= u7_t[64];
    u7_o[65] <= u7_t[65];
    u7_o[66] <= u7_t[66];
    u7_o[67] <= u7_t[67];
    u7_o[68] <= u7_t[68];
    u7_o[69] <= u7_t[69];
    u7_o[70] <= u7_t[70];
    u7_o[71] <= u7_t[71];
    u7_o[72] <= u7_t[72];
    u7_o[73] <= u7_t[73];
    u7_o[74] <= u7_t[74];
    u7_o[75] <= u7_t[75];
    u7_o[76] <= u7_t[76];
    u7_o[77] <= u7_t[77];
    u7_o[78] <= u7_t[78];
    u7_o[79] <= u7_t[79];
    u7_o[80] <= u7_t[80];
    u7_o[81] <= u7_t[81];
    u7_o[82] <= u7_t[82];
    u7_o[83] <= u7_t[83];
    u7_o[84] <= u7_t[84];
    u7_o[85] <= u7_t[85];
    u7_o[86] <= u7_t[86];
    u7_o[87] <= u7_t[87];
    u7_o[88] <= u7_t[88];
    u7_o[89] <= u7_t[89];
    u7_o[90] <= u7_t[90];
    u7_o[91] <= u7_t[91];
    u7_o[92] <= u7_t[92];
    u7_o[93] <= u7_t[93];
    u7_o[94] <= u7_t[94];
    u7_o[95] <= u7_t[95];
    u7_o[96] <= u7_t[96];
    u7_o[97] <= u7_t[97];
    u7_o[98] <= u7_t[98];
    u7_o[99] <= u7_t[99];
    u7_o[100] <= u7_t[100];
    u7_o[101] <= u7_t[101];
    u7_o[102] <= u7_t[102];
    u7_o[103] <= u7_t[103];
    u7_o[104] <= u7_t[104];
    u7_o[105] <= u7_t[105];
    u7_o[106] <= u7_t[106];
    u7_o[107] <= u7_t[107];
    u7_o[108] <= u7_t[108];
    u7_o[109] <= u7_t[109];
    u7_o[110] <= u7_t[110];
    u7_o[111] <= u7_t[111];
    u7_o[112] <= u7_t[112];
    u7_o[113] <= u7_t[113];
    u7_o[114] <= u7_t[114];
    u7_o[115] <= u7_t[115];
    u7_o[116] <= u7_t[116];
    u7_o[117] <= u7_t[117];
    u7_o[118] <= u7_t[118];
    u7_o[119] <= u7_t[119];
    u7_o[120] <= u7_t[120];
    u7_o[121] <= u7_t[121];
    u7_o[122] <= u7_t[122];
    u7_o[123] <= u7_t[123];
    u7_o[124] <= u7_t[124];
    u7_o[125] <= u7_t[125];
    u7_o[126] <= u7_t[126];
    u7_o[127] <= u7_t[127];
    u7_o[128] <= u7_t[128];
    u7_o[129] <= u7_t[129];
    u7_o[130] <= u7_t[130];
    u7_o[131] <= u7_t[131];
    u7_o[132] <= u7_t[132];
    u7_o[133] <= u7_t[133];
    u7_o[134] <= u7_t[134];
    u7_o[135] <= u7_t[135];
    u7_o[136] <= u7_t[136];
    u7_o[137] <= u7_t[137];
    u7_o[138] <= u7_t[138];
    u7_o[139] <= u7_t[139];
    u7_o[140] <= u7_t[140];
    u7_o[141] <= u7_t[141];
    u7_o[142] <= u7_t[142];
    u7_o[143] <= u7_t[143];
    u7_o[144] <= u7_t[144];
    u7_o[145] <= u7_t[145];
    u7_o[146] <= u7_t[146];
    u7_o[147] <= u7_t[147];
    u7_o[148] <= u7_t[148];
    u7_o[149] <= u7_t[149];
    u7_o[150] <= u7_t[150];
    u7_o[151] <= u7_t[151];
    u7_o[152] <= u7_t[152];
    u7_o[153] <= u7_t[153];
    u7_o[154] <= u7_t[154];
    u7_o[155] <= u7_t[155];
    u7_o[156] <= u7_t[156];
    u7_o[157] <= u7_t[157];
    u7_o[158] <= u7_t[158];
    u7_o[159] <= u7_t[159];
    u7_o[160] <= u7_t[160];
    u7_o[161] <= u7_t[161];
    u7_o[162] <= u7_t[162];
    u7_o[163] <= u7_t[163];
    u7_o[164] <= u7_t[164];
    u7_o[165] <= u7_t[165];
    u7_o[166] <= u7_t[166];
    u7_o[167] <= u7_t[167];
    u7_o[168] <= u7_t[168];
    u7_o[169] <= u7_t[169];
    u7_o[170] <= u7_t[170];
    u7_o[171] <= u7_t[171];
    u7_o[172] <= u7_t[172];
    u7_o[173] <= u7_t[173];
    u7_o[174] <= u7_t[174];
    u7_o[175] <= u7_t[175];
    u7_o[176] <= u7_t[176];
    u7_o[177] <= u7_t[177];
    u7_o[178] <= u7_t[178];
    u7_o[179] <= u7_t[179];
    u7_o[180] <= u7_t[180];
    u7_o[181] <= u7_t[181];
    u7_o[182] <= u7_t[182];
    u7_o[183] <= u7_t[183];
    u7_o[184] <= u7_t[184];
    u7_o[185] <= u7_t[185];
    u7_o[186] <= u7_t[186];
    u7_o[187] <= u7_t[187];
    u7_o[188] <= u7_t[188];
    u7_o[189] <= u7_t[189];
    u7_o[190] <= u7_t[190];
    u7_o[191] <= u7_t[191];
    u7_o[192] <= u7_t[192];
    u7_o[193] <= u7_t[193];
    u7_o[194] <= u7_t[194];
    u7_o[195] <= u7_t[195];
    u7_o[196] <= u7_t[196];
    u7_o[197] <= u7_t[197];
    u7_o[198] <= u7_t[198];
    u7_o[199] <= u7_t[199];
    u7_o[200] <= u7_t[200];
    u7_o[201] <= u7_t[201];
    u7_o[202] <= u7_t[202];
    u7_o[203] <= u7_t[203];
    u7_o[204] <= u7_t[204];
    u7_o[205] <= u7_t[205];
    u7_o[206] <= u7_t[206];
    u7_o[207] <= u7_t[207];
    u7_o[208] <= u7_t[208];
    u7_o[209] <= u7_t[209];
    u7_o[210] <= u7_t[210];
    u7_o[211] <= u7_t[211];
    u7_o[212] <= u7_t[212];
    u7_o[213] <= u7_t[213];
    u7_o[214] <= u7_t[214];
    u7_o[215] <= u7_t[215];
    u7_o[216] <= u7_t[216];
    u7_o[217] <= u7_t[217];
    u7_o[218] <= u7_t[218];
    u7_o[219] <= u7_t[219];
    u7_o[220] <= u7_t[220];
    u7_o[221] <= u7_t[221];
    u7_o[222] <= u7_t[222];
    u7_o[223] <= u7_t[223];
    u7_o[224] <= u7_t[224];
    u7_o[225] <= u7_t[225];
    u7_o[226] <= u7_t[226];
    u7_o[227] <= u7_t[227];
    u7_o[228] <= u7_t[228];
    u7_o[229] <= u7_t[229];
    u7_o[230] <= u7_t[230];
    u7_o[231] <= u7_t[231];
    u7_o[232] <= u7_t[232];
    u7_o[233] <= u7_t[233];
    u7_o[234] <= u7_t[234];
    u7_o[235] <= u7_t[235];
    u7_o[236] <= u7_t[236];
    u7_o[237] <= u7_t[237];
    u7_o[238] <= u7_t[238];
    u7_o[239] <= u7_t[239];
    u7_o[240] <= u7_t[240];
    u7_o[241] <= u7_t[241];
    u7_o[242] <= u7_t[242];
    u7_o[243] <= u7_t[243];
    u7_o[244] <= u7_t[244];
    u7_o[245] <= u7_t[245];
    u7_o[246] <= u7_t[246];
    u7_o[247] <= u7_t[247];
    u7_o[248] <= u7_t[248];
    u7_o[249] <= u7_t[249];
    u7_o[250] <= u7_t[250];
    u7_o[251] <= u7_t[251];
    u7_o[252] <= u7_t[252];
    u7_o[253] <= u7_t[253];
    u7_o[254] <= u7_t[254];
    u7_o[255] <= u7_t[255];
  end
  
  always@(*)begin
    for(i=0;i<510;i=i+1)begin
      if(i[0]==1'b0) u0_t[i] = u[i] ^ u[i+1];
      else           u0_t[i] = u[i];
    end
  end
  
  always@(*)begin
    for(i=0;i<508;i=i+1)begin
      if(i[1:0]<=2'd1) u1_t[i] = u0_t[i] ^ u0_t[i+2];
      else           u1_t[i] = u0_t[i];
    end
  end
  
  always@(*)begin
    for(i=0;i<504;i=i+1)begin
      if(i[2:0]<=3'd3) u2_t[i] = u1_t[i] ^ u1_t[i+4];
      else           u2_t[i] = u1_t[i];
    end
  end
  
  always@(*)begin
    for(i=0;i<496;i=i+1)begin
      if(i[3:0]<=4'd7) u3_t[i] = u2_t[i] ^ u2_t[i+8];
      else           u3_t[i] = u2_t[i];
    end
  end
  
  always@(*)begin
    for(i=0;i<480;i=i+1)begin
      if(i[4:0]<=5'd15) u4_t[i] = u3_t[i] ^ u3_t[i+16];
      else           u4_t[i] = u3_t[i];
    end
  end
  
  always@(*)begin
  /*
    for(i=0;i<512;i=i+1)begin
      if(i[5:0]<=6'd31) u5_t[i] = u4_t[i] ^ u4_t[i+32];
      else           u5_t[i] = u4_t[i];
    end
  */
    for(i=0;i<448;i=i+1)begin
      if(i[5:0]<=6'd31) u5_t[i] = u4_t[i] ^ u4_t[i+32];
      else           u5_t[i] = u4_t[i];
    end
  end
  
  always@(*)begin
  /*
    for(i=0;i<512;i=i+1)begin
      if(i[6:0]<=7'd63) u6_t[i] = u5_t[i] ^ u5_t[i+64];
      else           u6_t[i] = u5_t[i];
    end
  */
    for(i=0;i<384;i=i+1)begin
      if(i[6:0]<=7'd63) u6_t[i] = u5_t[i] ^ u5_t[i+64];
      else           u6_t[i] = u5_t[i];
    end
  end
  
  always@(*)begin
  /*
    for(i=0;i<512;i=i+1)begin
      if(i[7:0]<=8'd127) u7_t[i] = u6_t[i] ^ u6_t[i+128];
      else           u7_t[i] = u6_t[i];
    end
  */
    for(i=0;i<256;i=i+1)begin
      if(i[7:0]<=8'd127) u7_t[i] = u6_t[i] ^ u6_t[i+128];
      else           u7_t[i] = u6_t[i];
    end
  end
  
endmodule